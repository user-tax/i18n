       )Q���VmV;u�����ͽ8B�	
L| �z   
    ce'� �Pu	vbg{l��$��a!�Lu�=S9X�b]   
<p><a href="https://&lt;br host&gt;"><br host></a><br action>verifierings kod:<br code>.</p>    �u��ئ�&P��Xql�����ئU��zP9�ָ�=   
<p>Denna verifieringskod upphör att gälla om en timme.</p>    �m��l�J]�ɞt|w3�t3.����сa���&@   
<p>Om du inte har ansökt, ignorera detta e-postmeddelande.</p>    �>�������v��c�b�����1_Ǣ��_�����7   <p>[<br host>]<br action>verifierings kod:<br code></p>